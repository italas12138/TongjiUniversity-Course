
module selector_tb;
    reg [3:0] iC0,iC1,iC2,iC3;
    reg iS1,iS0;
    wire [3:0] oZ;
    selector41 uut(.iS0(iS0),.iS1(iS1),.iC0(iC0),.iC1(iC1),.iC2(iC2),.iC3(iC3),.oZ(oZ));
    initial
    begin
    iS1=0;
    iS0=0;
    iC0=4'b0000;
    iC1=4'b0000;
    iC2=4'b0000;
    iC3=4'b0000;
    #5;
    iC0=4'b1111;
    iC1=4'b0111;
    iC2=4'b0011;
    iC3=4'b0001;
    #5;
    iC0=4'b1111;
    iC1=4'b0000;
    iC2=4'b0000;
    iC3=4'b0000;
    #5;
    iC0=4'b0011;
    iC1=4'b0000;
    iC2=4'b0000;
    iC3=4'b0000;
     #5;
     iS0=1;
     iC0=4'b1111;
     iC1=4'b0111;
     iC2=4'b0011;
     iC3=4'b0001;
     #5;
     iC0=4'b0000;
     iC1=4'b0111;
     iC2=4'b0000;
     iC3=4'b0000;
     #5;
     iC0=4'b0000;
     iC1=4'b1111;
     iC2=4'b0000;
     iC3=4'b0000;
     #5;
     iS1=1;
     iS0=0;
     iC0=4'b1111;
     iC1=4'b0111;
     iC2=4'b0011;
     iC3=4'b0001;
     #5;
     iC0=4'b0000;
     iC1=4'b0000;
     iC2=4'b0011;
     iC3=4'b0000;
     #5;
     iC0=4'b0000;
     iC1=4'b0000;
     iC2=4'b1111;
     iC3=4'b0000;
     #5;
     iS0=1;
     iC0=4'b1111;
     iC1=4'b0111;
     iC2=4'b0011;
     iC3=4'b0001;
     #5;
     iC0=4'b0000;
     iC1=4'b0000;
     iC2=4'b0000;
     iC3=4'b0001;
     #5;
     iC0=4'b0000;
     iC1=4'b0000;
     iC2=4'b0000;
     iC3=4'b1111;
     end
endmodule
